netcdf basic {
dimensions:
}
